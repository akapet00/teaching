* C:\Users\Maja-FESB\Documents\Schematicpreslusavanje.sch

* Schematics Version 9.1 - Web Update 1
* Tue Dec 19 12:41:55 2017



** Analysis setup **
.ac DEC 101 10 10000.00K


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematicpreslusavanje.net"
.INC "Schematicpreslusavanje.als"


.probe


.END
