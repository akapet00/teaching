* C:\Users\Maja-FESB\Documents\Schematic2.sch

* Schematics Version 9.1 - Web Update 1
* Fri Jan 18 09:13:47 2019



** Analysis setup **
.ac DEC 101 10 100.00K


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic2.net"
.INC "Schematic2.als"


.probe


.END
