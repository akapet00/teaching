* C:\Users\Maja-FESB\Documents\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Thu Dec 06 16:08:23 2018



** Analysis setup **
.tran 0s 500e-6s 0 100ns


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
