* C:\Users\Maja-FESB\Documents\Schematic3.sch

* Schematics Version 9.1 - Web Update 1
* Thu Jan 17 16:02:22 2019



** Analysis setup **
.tran 0 500e-6 0 100ns


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic3.net"
.INC "Schematic3.als"


.probe


.END
