* C:\Users\Maja-FESB\Documents\Schematictl.sch

* Schematics Version 9.1 - Web Update 1
* Tue Dec 19 14:12:29 2017



** Analysis setup **
.tran 0s 500e-6s 0 100ns


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematictl.net"
.INC "Schematictl.als"


.probe


.END
